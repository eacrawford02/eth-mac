// Copyright (C) 2023 Ewen Crawford

module tb();
  tb_afifo afifo_test();
endmodule
